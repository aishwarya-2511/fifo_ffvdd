`include "Sync_FIFO.v"
`include "fifo_trans.sv"
`include "fifo_gen.sv"
`include "fifo_intf.sv"
`include "fifo_bfm.sv"
`include "fifo_env.sv"
`include "fifo_test.sv"
`include "fifo_top.sv"





